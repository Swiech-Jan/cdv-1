<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>2.41875,0.2875,52.0313,-33.7438</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>9,-11</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>9,-14.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>9,-21</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>18,-2.5</position>
<gparam>LABEL_TEXT Y = !ABD + A!D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>5,-10.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>5,-14</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>5.5,-20.5</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_AND3</type>
<position>26.5,-13.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>7 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>27,-24.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AE_OR2</type>
<position>35.5,-18</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>43.5,-17</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_INVERTER</type>
<position>18.5,-11.5</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_INVERTER</type>
<position>18,-26</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-17,31,-13.5</points>
<intersection>-17 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-17,32.5,-17</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-13.5,31,-13.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-24.5,31,-19</points>
<intersection>-24.5 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-19,32.5,-19</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-24.5,31,-24.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,-18,40.5,-18</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-11.5,13,-11</points>
<intersection>-11.5 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-11.5,15.5,-11.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection>
<intersection>14.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-11,13,-11</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>13 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14.5,-23.5,14.5,-11.5</points>
<intersection>-23.5 4</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>14.5,-23.5,24,-23.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>14.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-11.5,23.5,-11.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-14.5,17,-13.5</points>
<intersection>-14.5 2</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-13.5,23.5,-13.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-14.5,17,-14.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-21,17,-15.5</points>
<intersection>-21 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-15.5,23.5,-15.5</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-21,17,-21</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>13 3</intersection>
<intersection>17 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13,-26,13,-21</points>
<intersection>-26 4</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>13,-26,15,-26</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>13 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-26,22.5,-25.5</points>
<intersection>-26 2</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-25.5,24,-25.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-26,22.5,-26</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-2.475,1.45,63.675,-43.925</PageViewport>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>13.5,-3.5</position>
<gparam>LABEL_TEXT Y = !AB + !ACD</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>9.5,-11</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>9.5,-14.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>9.5,-18</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_TOGGLE</type>
<position>9.5,-21.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>6.5,-10.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>6.5,-14</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>6.5,-17.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>6.5,-21</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AE_OR2</type>
<position>43.5,-33.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>53.5,-32.5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_AND2</type>
<position>34.5,-28</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND3</type>
<position>34,-36.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>15 </input>
<input>
<ID>IN_2</ID>16 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_INVERTER</type>
<position>26.5,-25.5</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-33.5,50.5,-33.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-32.5,39,-28</points>
<intersection>-32.5 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-32.5,40.5,-32.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-28,39,-28</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-36.5,38.5,-34.5</points>
<intersection>-36.5 2</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-34.5,40.5,-34.5</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,-36.5,38.5,-36.5</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>7</ID>
<points>30,-34.5,30,-25.5</points>
<intersection>-34.5 8</intersection>
<intersection>-27 9</intersection>
<intersection>-25.5 10</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>30,-34.5,31,-34.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>30 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>30,-27,31.5,-27</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>30 7</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>29.5,-25.5,30,-25.5</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>30 7</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-25.5,22,-11</points>
<intersection>-25.5 2</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,-11,22,-11</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-25.5,23.5,-25.5</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-29,21,-14.5</points>
<intersection>-29 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-29,31.5,-29</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-14.5,21,-14.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-36.5,19.5,-18</points>
<intersection>-36.5 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,-18,19.5,-18</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-36.5,31,-36.5</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-38.5,17.5,-21.5</points>
<intersection>-38.5 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,-21.5,17.5,-21.5</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-38.5,31,-38.5</points>
<connection>
<GID>44</GID>
<name>IN_2</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-2.475,1.45,63.675,-43.925</PageViewport>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>15.5,-3</position>
<gparam>LABEL_TEXT Y = !A (B+C)(B+D)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_AND3</type>
<position>40,-31.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>22 </input>
<input>
<ID>IN_2</ID>24 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>52</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>50,-30.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>4.5,-8.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_TOGGLE</type>
<position>7.5,-9</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>4.5,-12</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_TOGGLE</type>
<position>7.5,-12.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>59</ID>
<type>AA_LABEL</type>
<position>4.5,-15.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_TOGGLE</type>
<position>7.5,-16</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>4.5,-19</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_TOGGLE</type>
<position>7.5,-19.5</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_INVERTER</type>
<position>26,-23</position>
<input>
<ID>IN_0</ID>19 </input>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>66</ID>
<type>AE_OR2</type>
<position>25.5,-31.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>68</ID>
<type>AE_OR2</type>
<position>25.5,-37.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-31.5,47,-31.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<connection>
<GID>50</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-29.5,37,-29.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>29 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>29,-29.5,29,-23</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>-29.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-23,18,-9</points>
<intersection>-23 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,-9,18,-9</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-23,23,-23</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-30.5,16,-12.5</points>
<intersection>-30.5 1</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-30.5,22.5,-30.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection>
<intersection>19 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-12.5,16,-12.5</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>16 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>19,-36.5,19,-30.5</points>
<intersection>-36.5 4</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-36.5,22.5,-36.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>19 3</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-32.5,14,-16</points>
<intersection>-32.5 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14,-32.5,22.5,-32.5</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-16,14,-16</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-31.5,37,-31.5</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<connection>
<GID>50</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-38.5,12,-19.5</points>
<intersection>-38.5 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,-19.5,12,-19.5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-38.5,22.5,-38.5</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>12 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-37.5,32.5,-33.5</points>
<intersection>-37.5 2</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-33.5,37,-33.5</points>
<connection>
<GID>50</GID>
<name>IN_2</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-37.5,32.5,-37.5</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,0,88.2,-60.5</PageViewport>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>27,-2</position>
<gparam>LABEL_TEXT Uklad sumujacy (funkcja S oraz C)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>3,-10.5</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>11.5,-10.5</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_TOGGLE</type>
<position>21,-10.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>3,-7</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>AA_LABEL</type>
<position>12,-7</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>21,-7</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>AE_OR2</type>
<position>62,-30</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>72.5,-29</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_AND2</type>
<position>52.5,-27</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>87</ID>
<type>AA_AND2</type>
<position>52.5,-34</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>AO_XNOR2</type>
<position>32,-21.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>91</ID>
<type>AA_INVERTER</type>
<position>43.5,-36</position>
<input>
<ID>IN_0</ID>29 </input>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>93</ID>
<type>AI_XOR2</type>
<position>32,-33</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>72.5,-22</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AE_OR3</type>
<position>48.5,-48.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>39 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_AND2</type>
<position>34,-42</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>100</ID>
<type>AA_AND2</type>
<position>34,-48.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_AND2</type>
<position>34,-55</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>103</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>72.5,-47.5</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>72.5,-41</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65,-30,69.5,-30</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<connection>
<GID>84</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-29,57,-27</points>
<intersection>-29 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57,-29,59,-29</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-27,57,-27</points>
<connection>
<GID>86</GID>
<name>OUT</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-34,57,-31</points>
<intersection>-34 2</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57,-31,59,-31</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-34,57,-34</points>
<connection>
<GID>87</GID>
<name>OUT</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-26,36.5,-21.5</points>
<intersection>-26 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-26,49.5,-26</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-21.5,36.5,-21.5</points>
<connection>
<GID>89</GID>
<name>OUT</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-28,24.5,-10.5</points>
<intersection>-28 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-10.5,24.5,-10.5</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-28,49.5,-28</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection>
<intersection>26.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>26.5,-43,26.5,-28</points>
<intersection>-43 5</intersection>
<intersection>-36 4</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>26.5,-36,40.5,-36</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>26.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>26.5,-43,31,-43</points>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<intersection>26.5 3</intersection>
<intersection>29.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>29.5,-56,29.5,-43</points>
<intersection>-56 7</intersection>
<intersection>-43 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>29.5,-56,31,-56</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>29.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-20.5,7.5,-10.5</points>
<intersection>-20.5 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-10.5,7.5,-10.5</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>7.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7.5,-20.5,29,-20.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>7.5 0</intersection>
<intersection>10.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>10.5,-32,10.5,-20.5</points>
<intersection>-32 4</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>10.5,-32,29,-32</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>10.5 3</intersection>
<intersection>14 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>14,-41,14,-32</points>
<intersection>-41 6</intersection>
<intersection>-32 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>14,-41,31,-41</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>14 5</intersection>
<intersection>17.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>17.5,-47.5,17.5,-41</points>
<intersection>-47.5 8</intersection>
<intersection>-41 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>17.5,-47.5,31,-47.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>17.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-22.5,16.5,-10.5</points>
<intersection>-22.5 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13.5,-10.5,16.5,-10.5</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-22.5,29,-22.5</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<intersection>16.5 0</intersection>
<intersection>19.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>19.5,-34,19.5,-22.5</points>
<intersection>-34 4</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19.5,-34,29,-34</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<intersection>19.5 3</intersection>
<intersection>22 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>22,-49.5,22,-34</points>
<intersection>-49.5 6</intersection>
<intersection>-34 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>22,-49.5,31,-49.5</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>22 5</intersection>
<intersection>25 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>25,-54,25,-49.5</points>
<intersection>-54 8</intersection>
<intersection>-49.5 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>25,-54,31,-54</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>25 7</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-36,49.5,-36</points>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection>
<intersection>49.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>49.5,-36,49.5,-35</points>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<intersection>-36 1</intersection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-33,49.5,-33</points>
<connection>
<GID>93</GID>
<name>OUT</name></connection>
<connection>
<GID>87</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,-48.5,69.5,-48.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<connection>
<GID>97</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-46.5,41,-42</points>
<intersection>-46.5 1</intersection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-46.5,45.5,-46.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,-42,41,-42</points>
<connection>
<GID>99</GID>
<name>OUT</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-48.5,45.5,-48.5</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<connection>
<GID>100</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-55,41,-50.5</points>
<intersection>-55 2</intersection>
<intersection>-50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-50.5,45.5,-50.5</points>
<connection>
<GID>97</GID>
<name>IN_2</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,-55,41,-55</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>0,0,88.2,-60.5</PageViewport>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>9.5,-2</position>
<gparam>LABEL_TEXT Polsumator</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AA_TOGGLE</type>
<position>6,-6.5</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_LABEL</type>
<position>3,-6</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>AA_TOGGLE</type>
<position>6,-10.5</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>3,-10</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>AE_OR2</type>
<position>41.5,-18.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_AND2</type>
<position>41,-34.5</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>54,-14.5</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>119</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>53.5,-33.5</position>
<input>
<ID>IN_0</ID>46 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>120</ID>
<type>AA_LABEL</type>
<position>43.5,-11</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>121</ID>
<type>AA_LABEL</type>
<position>43.5,-30.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>AA_AND2</type>
<position>28,-14</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_AND2</type>
<position>28,-27.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_INVERTER</type>
<position>16.5,-17</position>
<input>
<ID>IN_0</ID>44 </input>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_INVERTER</type>
<position>18,-24</position>
<input>
<ID>IN_0</ID>40 </input>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-33.5,12,-6.5</points>
<intersection>-33.5 5</intersection>
<intersection>-24 3</intersection>
<intersection>-13 1</intersection>
<intersection>-6.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-13,25,-13</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-6.5,12,-6.5</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>12,-24,15,-24</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>12,-33.5,38,-33.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>12 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-17.5,34.5,-14</points>
<intersection>-17.5 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-17.5,38.5,-17.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-14,34.5,-14</points>
<connection>
<GID>124</GID>
<name>OUT</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-27.5,35,-19.5</points>
<intersection>-27.5 3</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-19.5,38.5,-19.5</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31,-27.5,35,-27.5</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-17,22,-15</points>
<intersection>-17 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-15,25,-15</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-17,22,-17</points>
<connection>
<GID>127</GID>
<name>OUT_0</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,-17,8.5,-10.5</points>
<intersection>-17 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,-10.5,8.5,-10.5</points>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-17,13.5,-17</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>8.5 0</intersection>
<intersection>10 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>10,-28.5,10,-17</points>
<intersection>-28.5 4</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>10,-28.5,25,-28.5</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>10 3</intersection>
<intersection>17 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>17,-35.5,17,-28.5</points>
<intersection>-35.5 6</intersection>
<intersection>-28.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>17,-35.5,38,-35.5</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>17 5</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21,-24,25,-24</points>
<connection>
<GID>128</GID>
<name>OUT_0</name></connection>
<intersection>25 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>25,-26.5,25,-24</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>-24 1</intersection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-34.5,50.5,-34.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<connection>
<GID>116</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-18.5,47.5,-15.5</points>
<intersection>-18.5 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-15.5,51,-15.5</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>44.5,-18.5,47.5,-18.5</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>-2.475,1.45,63.675,-43.925</PageViewport>
<gate>
<ID>130</ID>
<type>AA_LABEL</type>
<position>4.5,-5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AA_TOGGLE</type>
<position>8,-5.5</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_LABEL</type>
<position>10,-1.5</position>
<gparam>LABEL_TEXT Polsumator</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>AA_LABEL</type>
<position>4.5,-9</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>AA_TOGGLE</type>
<position>8,-9.5</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>138</ID>
<type>AI_XOR2</type>
<position>21,-15</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>140</ID>
<type>AA_AND2</type>
<position>20.5,-24</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>29.5,-14</position>
<input>
<ID>IN_0</ID>50 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>143</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>29.5,-23</position>
<input>
<ID>IN_0</ID>51 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_LABEL</type>
<position>29.5,-7.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>145</ID>
<type>AA_LABEL</type>
<position>29.5,-27.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-14,14.5,-5.5</points>
<intersection>-14 1</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-14,18,-14</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection>
<intersection>16 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10,-5.5,14.5,-5.5</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16,-23,16,-14</points>
<intersection>-23 4</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>16,-23,17.5,-23</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>16 3</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-16,12,-9.5</points>
<intersection>-16 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-16,18,-16</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>12 0</intersection>
<intersection>14.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10,-9.5,12,-9.5</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<intersection>12 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14.5,-25,14.5,-16</points>
<intersection>-25 4</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>14.5,-25,17.5,-25</points>
<connection>
<GID>140</GID>
<name>IN_1</name></connection>
<intersection>14.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-15,26.5,-15</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23.5,-24,26.5,-24</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<connection>
<GID>140</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>0,0,88.2,-60.5</PageViewport>
<gate>
<ID>147</ID>
<type>AA_LABEL</type>
<position>7.5,-2</position>
<gparam>LABEL_TEXT Sumator</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>AA_AND3</type>
<position>12,-10.5</position>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_LABEL</type>
<position>7.5,-8</position>
<gparam>LABEL_TEXT !A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>153</ID>
<type>AA_LABEL</type>
<position>7.5,-10</position>
<gparam>LABEL_TEXT !B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>AA_LABEL</type>
<position>6.5,-12</position>
<gparam>LABEL_TEXT C (IN)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>AA_AND3</type>
<position>12,-20</position>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>156</ID>
<type>AA_LABEL</type>
<position>7.5,-17.5</position>
<gparam>LABEL_TEXT !A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>AA_LABEL</type>
<position>7.5,-19.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>AA_LABEL</type>
<position>6.5,-21.5</position>
<gparam>LABEL_TEXT !C (IN)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>AA_AND3</type>
<position>12,-28.5</position>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>160</ID>
<type>AA_LABEL</type>
<position>7.5,-26</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>AA_LABEL</type>
<position>7.5,-28</position>
<gparam>LABEL_TEXT !B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>AA_LABEL</type>
<position>6.5,-30</position>
<gparam>LABEL_TEXT !C (IN)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>AA_AND3</type>
<position>12,-37</position>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>164</ID>
<type>AA_LABEL</type>
<position>7.5,-34.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>AA_LABEL</type>
<position>7.5,-36.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>AA_LABEL</type>
<position>6.5,-38.5</position>
<gparam>LABEL_TEXT C (IN)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AE_OR4</type>
<position>31.5,-22</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>55 </input>
<input>
<ID>IN_2</ID>56 </input>
<input>
<ID>IN_3</ID>57 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_LABEL</type>
<position>36.5,-21.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>AA_AND2</type>
<position>50.5,-16</position>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_LABEL</type>
<position>46,-14.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>177</ID>
<type>AA_LABEL</type>
<position>46,-16.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>AA_AND2</type>
<position>50.5,-23</position>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_LABEL</type>
<position>46,-21.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>AA_LABEL</type>
<position>46,-23.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>181</ID>
<type>AA_AND2</type>
<position>50.5,-30</position>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>182</ID>
<type>AA_LABEL</type>
<position>46,-28.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>AA_LABEL</type>
<position>46,-30.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>185</ID>
<type>AE_OR3</type>
<position>64,-23</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>59 </input>
<input>
<ID>IN_2</ID>60 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>70.5,-22.5</position>
<gparam>LABEL_TEXT C (OUT)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-19,21.5,-10.5</points>
<intersection>-19 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-10.5,21.5,-10.5</points>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-19,28.5,-19</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-21,21.5,-20</points>
<intersection>-21 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-20,21.5,-20</points>
<connection>
<GID>155</GID>
<name>OUT</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-21,28.5,-21</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-28.5,21.5,-23</points>
<intersection>-28.5 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-28.5,21.5,-28.5</points>
<connection>
<GID>159</GID>
<name>OUT</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-23,28.5,-23</points>
<connection>
<GID>170</GID>
<name>IN_2</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-37,23.5,-25</points>
<intersection>-37 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-37,23.5,-37</points>
<connection>
<GID>163</GID>
<name>OUT</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23.5,-25,28.5,-25</points>
<connection>
<GID>170</GID>
<name>IN_3</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-21,57,-16</points>
<intersection>-21 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57,-21,61,-21</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53.5,-16,57,-16</points>
<connection>
<GID>174</GID>
<name>OUT</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-23,61,-23</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<connection>
<GID>178</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-30,57,-25</points>
<intersection>-30 2</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57,-25,61,-25</points>
<connection>
<GID>185</GID>
<name>IN_2</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53.5,-30,57,-30</points>
<connection>
<GID>181</GID>
<name>OUT</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire></page 6>
<page 7>
<PageViewport>0,0,88.2,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,88.2,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,88.2,-60.5</PageViewport></page 9></circuit>