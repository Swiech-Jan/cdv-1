<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-0.100358,6.95439,316.759,-156.643</PageViewport>
<gate>
<ID>8</ID>
<type>DD_KEYPAD_HEX</type>
<position>46,-69</position>
<output>
<ID>OUT_0</ID>3 </output>
<output>
<ID>OUT_1</ID>4 </output>
<output>
<ID>OUT_2</ID>5 </output>
<output>
<ID>OUT_3</ID>6 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>62,-78</position>
<input>
<ID>N_in3</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>59,-78</position>
<input>
<ID>N_in3</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>56,-78</position>
<input>
<ID>N_in3</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>53,-78</position>
<input>
<ID>N_in3</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AI_XOR2</type>
<position>79,-36.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_AND2</type>
<position>74,-36.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>AE_OR2</type>
<position>75,-24</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>AI_XOR2</type>
<position>85,-30</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_AND2</type>
<position>80,-30</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>90</ID>
<type>HA_JUNC_2</type>
<position>73,-44</position>
<input>
<ID>N_in0</ID>85 </input>
<input>
<ID>N_in1</ID>43 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>91</ID>
<type>HA_JUNC_2</type>
<position>80,-44</position>
<input>
<ID>N_in0</ID>4 </input>
<input>
<ID>N_in1</ID>42 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>92</ID>
<type>HA_JUNC_2</type>
<position>86,-44</position>
<input>
<ID>N_in0</ID>65 </input>
<input>
<ID>N_in1</ID>46 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>94</ID>
<type>AA_LABEL</type>
<position>88.5,-43.5</position>
<gparam>LABEL_TEXT CIN</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>81.5,-43.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>74.5,-43.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>98</ID>
<type>HA_JUNC_2</type>
<position>75,-20</position>
<input>
<ID>N_in0</ID>50 </input>
<input>
<ID>N_in1</ID>83 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>0,0</position>
<gparam>LABEL_TEXT CIN</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>101</ID>
<type>HA_JUNC_2</type>
<position>85,-20</position>
<input>
<ID>N_in0</ID>53 </input>
<input>
<ID>N_in1</ID>89 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>86.5,-19.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>103</ID>
<type>AA_LABEL</type>
<position>78,-19.5</position>
<gparam>LABEL_TEXT COUT</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>108</ID>
<type>AI_XOR2</type>
<position>103,-36.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_AND2</type>
<position>98,-36.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>HA_JUNC_2</type>
<position>97,-44</position>
<input>
<ID>N_in0</ID>84 </input>
<input>
<ID>N_in1</ID>58 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>114</ID>
<type>HA_JUNC_2</type>
<position>104,-44</position>
<input>
<ID>N_in0</ID>3 </input>
<input>
<ID>N_in1</ID>57 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>117</ID>
<type>AA_LABEL</type>
<position>105.5,-43.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>98.5,-43.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>119</ID>
<type>HA_JUNC_2</type>
<position>98,-30</position>
<input>
<ID>N_in0</ID>2 </input>
<input>
<ID>N_in1</ID>65 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>120</ID>
<type>HA_JUNC_2</type>
<position>109,-30</position>
<input>
<ID>N_in0</ID>1 </input>
<input>
<ID>N_in1</ID>88 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>121</ID>
<type>AA_LABEL</type>
<position>110.5,-29.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>122</ID>
<type>AA_LABEL</type>
<position>101,-29.5</position>
<gparam>LABEL_TEXT COUT</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>123</ID>
<type>AI_XOR2</type>
<position>31,-36.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>124</ID>
<type>AA_AND2</type>
<position>26,-36.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>125</ID>
<type>AE_OR2</type>
<position>27,-24</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>71 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>AI_XOR2</type>
<position>37,-30</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_AND2</type>
<position>32,-30</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>128</ID>
<type>HA_JUNC_2</type>
<position>25,-44</position>
<input>
<ID>N_in0</ID>87 </input>
<input>
<ID>N_in1</ID>67 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>129</ID>
<type>HA_JUNC_2</type>
<position>32,-44</position>
<input>
<ID>N_in0</ID>6 </input>
<input>
<ID>N_in1</ID>66 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>130</ID>
<type>HA_JUNC_2</type>
<position>38,-44</position>
<input>
<ID>N_in0</ID>82 </input>
<input>
<ID>N_in1</ID>69 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>131</ID>
<type>AA_LABEL</type>
<position>40.5,-43.5</position>
<gparam>LABEL_TEXT CIN</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>132</ID>
<type>AA_LABEL</type>
<position>33.5,-43.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>133</ID>
<type>AA_LABEL</type>
<position>26.5,-43.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>134</ID>
<type>HA_JUNC_2</type>
<position>27,-20</position>
<input>
<ID>N_in0</ID>72 </input>
<input>
<ID>N_in1</ID>92 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>135</ID>
<type>HA_JUNC_2</type>
<position>37,-20</position>
<input>
<ID>N_in0</ID>73 </input>
<input>
<ID>N_in1</ID>91 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>136</ID>
<type>AA_LABEL</type>
<position>38.5,-19.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>137</ID>
<type>AA_LABEL</type>
<position>30,-19.5</position>
<gparam>LABEL_TEXT COUT</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>138</ID>
<type>AI_XOR2</type>
<position>55,-36.5</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>139</ID>
<type>AA_AND2</type>
<position>50,-36.5</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>140</ID>
<type>AE_OR2</type>
<position>51,-24</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>141</ID>
<type>AI_XOR2</type>
<position>61,-30</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>77 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_AND2</type>
<position>56,-30</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>77 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>143</ID>
<type>HA_JUNC_2</type>
<position>49,-44</position>
<input>
<ID>N_in0</ID>86 </input>
<input>
<ID>N_in1</ID>75 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>144</ID>
<type>HA_JUNC_2</type>
<position>56,-44</position>
<input>
<ID>N_in0</ID>5 </input>
<input>
<ID>N_in1</ID>74 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>145</ID>
<type>HA_JUNC_2</type>
<position>62,-44</position>
<input>
<ID>N_in0</ID>83 </input>
<input>
<ID>N_in1</ID>77 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>146</ID>
<type>AA_LABEL</type>
<position>64.5,-43.5</position>
<gparam>LABEL_TEXT CIN</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>147</ID>
<type>AA_LABEL</type>
<position>57.5,-43.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>148</ID>
<type>AA_LABEL</type>
<position>50.5,-43.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>149</ID>
<type>HA_JUNC_2</type>
<position>51,-20</position>
<input>
<ID>N_in0</ID>80 </input>
<input>
<ID>N_in1</ID>82 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>150</ID>
<type>HA_JUNC_2</type>
<position>61,-20</position>
<input>
<ID>N_in0</ID>81 </input>
<input>
<ID>N_in1</ID>90 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>151</ID>
<type>AA_LABEL</type>
<position>62.5,-19.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>152</ID>
<type>AA_LABEL</type>
<position>54,-19.5</position>
<gparam>LABEL_TEXT COUT</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>153</ID>
<type>DD_KEYPAD_HEX</type>
<position>81,-69</position>
<output>
<ID>OUT_0</ID>84 </output>
<output>
<ID>OUT_1</ID>85 </output>
<output>
<ID>OUT_2</ID>86 </output>
<output>
<ID>OUT_3</ID>87 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>154</ID>
<type>GA_LED</type>
<position>97,-78</position>
<input>
<ID>N_in3</ID>84 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>GA_LED</type>
<position>94,-78</position>
<input>
<ID>N_in3</ID>85 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>GA_LED</type>
<position>91,-78</position>
<input>
<ID>N_in3</ID>86 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>GA_LED</type>
<position>88,-78</position>
<input>
<ID>N_in3</ID>87 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>121.5,-14</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>89 </input>
<input>
<ID>IN_2</ID>90 </input>
<input>
<ID>IN_3</ID>91 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>160</ID>
<type>GA_LED</type>
<position>109,-8</position>
<input>
<ID>N_in2</ID>88 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>GA_LED</type>
<position>106,-8</position>
<input>
<ID>N_in0</ID>89 </input>
<input>
<ID>N_in2</ID>89 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>GA_LED</type>
<position>103,-8</position>
<input>
<ID>N_in2</ID>90 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>GA_LED</type>
<position>100,-8</position>
<input>
<ID>N_in2</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>GA_LED</type>
<position>95,-8</position>
<input>
<ID>N_in2</ID>92 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>169</ID>
<type>AA_LABEL</type>
<position>81,-76.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AA_LABEL</type>
<position>46,-76.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>AA_LABEL</type>
<position>62,-80</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>AA_LABEL</type>
<position>97,-80</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>AA_LABEL</type>
<position>59,-80</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>AA_LABEL</type>
<position>56,-80</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>AA_LABEL</type>
<position>53,-80</position>
<gparam>LABEL_TEXT 8</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>176</ID>
<type>AA_LABEL</type>
<position>94,-80</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>177</ID>
<type>AA_LABEL</type>
<position>91,-80</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>AA_LABEL</type>
<position>88,-80</position>
<gparam>LABEL_TEXT 8</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>179</ID>
<type>AA_LABEL</type>
<position>109,-5.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>AA_LABEL</type>
<position>106,-5.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>181</ID>
<type>AA_LABEL</type>
<position>103,-5.5</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>182</ID>
<type>AA_LABEL</type>
<position>100,-5.5</position>
<gparam>LABEL_TEXT 8</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>AA_LABEL</type>
<position>95,-5.5</position>
<gparam>LABEL_TEXT 16</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,-32,109,-31</points>
<connection>
<GID>120</GID>
<name>N_in0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>103,-33.5,103,-32</points>
<connection>
<GID>108</GID>
<name>OUT</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>103,-32,109,-32</points>
<intersection>103 1</intersection>
<intersection>109 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-33.5,98,-31</points>
<connection>
<GID>109</GID>
<name>OUT</name></connection>
<connection>
<GID>119</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51,-72,62,-72</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>62 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>62,-77,62,-53.5</points>
<connection>
<GID>10</GID>
<name>N_in3</name></connection>
<intersection>-72 1</intersection>
<intersection>-53.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>62,-53.5,104,-53.5</points>
<intersection>62 3</intersection>
<intersection>104 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>104,-53.5,104,-45</points>
<connection>
<GID>114</GID>
<name>N_in0</name></connection>
<intersection>-53.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-77,59,-51.5</points>
<connection>
<GID>12</GID>
<name>N_in3</name></connection>
<intersection>-70 1</intersection>
<intersection>-51.5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-70,59,-70</points>
<connection>
<GID>8</GID>
<name>OUT_1</name></connection>
<intersection>59 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>59,-51.5,80,-51.5</points>
<intersection>59 0</intersection>
<intersection>80 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>80,-51.5,80,-45</points>
<connection>
<GID>91</GID>
<name>N_in0</name></connection>
<intersection>-51.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-77,56,-45</points>
<connection>
<GID>144</GID>
<name>N_in0</name></connection>
<connection>
<GID>14</GID>
<name>N_in3</name></connection>
<intersection>-68 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>51,-68,56,-68</points>
<connection>
<GID>8</GID>
<name>OUT_2</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-77,53,-57.5</points>
<connection>
<GID>16</GID>
<name>N_in3</name></connection>
<intersection>-66 6</intersection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-57.5,53,-57.5</points>
<intersection>32 4</intersection>
<intersection>53 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>32,-57.5,32,-45</points>
<connection>
<GID>129</GID>
<name>N_in0</name></connection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>51,-66,53,-66</points>
<connection>
<GID>8</GID>
<name>OUT_3</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-43,80,-39.5</points>
<connection>
<GID>75</GID>
<name>IN_1</name></connection>
<connection>
<GID>91</GID>
<name>N_in1</name></connection>
<intersection>-40.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>75,-40.5,80,-40.5</points>
<intersection>75 5</intersection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>75,-40.5,75,-39.5</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>-40.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-42,78,-39.5</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>-42 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>73,-43,73,-39.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<connection>
<GID>90</GID>
<name>N_in1</name></connection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>73,-42,78,-42</points>
<intersection>73 1</intersection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>79,-33.5,84,-33.5</points>
<connection>
<GID>75</GID>
<name>OUT</name></connection>
<intersection>79 16</intersection>
<intersection>84 17</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>79,-33.5,79,-33</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>-33.5 3</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>84,-33.5,84,-33</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>-33.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-43,86,-33</points>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<connection>
<GID>92</GID>
<name>N_in1</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>81,-34.5,86,-34.5</points>
<intersection>81 4</intersection>
<intersection>86 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>81,-34.5,81,-33</points>
<connection>
<GID>84</GID>
<name>IN_1</name></connection>
<intersection>-34.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-33.5,74,-27</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<connection>
<GID>82</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>76,-27,80,-27</points>
<connection>
<GID>84</GID>
<name>OUT</name></connection>
<connection>
<GID>82</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-21,75,-21</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<connection>
<GID>98</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-27,85,-21</points>
<connection>
<GID>83</GID>
<name>OUT</name></connection>
<connection>
<GID>101</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-43,104,-39.5</points>
<connection>
<GID>114</GID>
<name>N_in1</name></connection>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>-40 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>99,-40,104,-40</points>
<intersection>99 5</intersection>
<intersection>104 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>99,-40,99,-39.5</points>
<connection>
<GID>109</GID>
<name>IN_1</name></connection>
<intersection>-40 4</intersection></vsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-42,102,-39.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-42 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>97,-43,97,-39.5</points>
<connection>
<GID>113</GID>
<name>N_in1</name></connection>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97,-42,102,-42</points>
<intersection>97 1</intersection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-46,92.5,-27</points>
<intersection>-46 2</intersection>
<intersection>-27 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>86,-46,86,-45</points>
<connection>
<GID>92</GID>
<name>N_in0</name></connection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>86,-46,92.5,-46</points>
<intersection>86 1</intersection>
<intersection>92.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>92.5,-27,98,-27</points>
<intersection>92.5 0</intersection>
<intersection>98 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>98,-29,98,-27</points>
<connection>
<GID>119</GID>
<name>N_in1</name></connection>
<intersection>-27 3</intersection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-43,32,-39.5</points>
<connection>
<GID>129</GID>
<name>N_in1</name></connection>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<intersection>-40.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>27,-40.5,32,-40.5</points>
<intersection>27 5</intersection>
<intersection>32 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>27,-40.5,27,-39.5</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>-40.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-42,30,-39.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>-42 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>25,-43,25,-39.5</points>
<connection>
<GID>128</GID>
<name>N_in1</name></connection>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>25,-42,30,-42</points>
<intersection>25 1</intersection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>31,-33.5,36,-33.5</points>
<connection>
<GID>123</GID>
<name>OUT</name></connection>
<intersection>31 16</intersection>
<intersection>36 17</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>31,-33.5,31,-33</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>-33.5 3</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>36,-33.5,36,-33</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>-33.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-43,38,-33</points>
<connection>
<GID>130</GID>
<name>N_in1</name></connection>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>33,-34.5,38,-34.5</points>
<intersection>33 4</intersection>
<intersection>38 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>33,-34.5,33,-33</points>
<connection>
<GID>127</GID>
<name>IN_1</name></connection>
<intersection>-34.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-33.5,26,-27</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<connection>
<GID>124</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>28,-27,32,-27</points>
<connection>
<GID>127</GID>
<name>OUT</name></connection>
<connection>
<GID>125</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-21,27,-21</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<connection>
<GID>134</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-27,37,-21</points>
<connection>
<GID>135</GID>
<name>N_in0</name></connection>
<connection>
<GID>126</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-43,56,-39.5</points>
<connection>
<GID>144</GID>
<name>N_in1</name></connection>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>-40 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>51,-40,56,-40</points>
<intersection>51 5</intersection>
<intersection>56 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>51,-40,51,-39.5</points>
<connection>
<GID>139</GID>
<name>IN_1</name></connection>
<intersection>-40 4</intersection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-42,54,-39.5</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>-42 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>49,-43,49,-39.5</points>
<connection>
<GID>143</GID>
<name>N_in1</name></connection>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>49,-42,54,-42</points>
<intersection>49 1</intersection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>55,-33.5,60,-33.5</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<intersection>55 16</intersection>
<intersection>60 17</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>55,-33.5,55,-33</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>-33.5 3</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>60,-33.5,60,-33</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>-33.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-43,62,-33</points>
<connection>
<GID>145</GID>
<name>N_in1</name></connection>
<connection>
<GID>141</GID>
<name>IN_1</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>57,-34.5,62,-34.5</points>
<intersection>57 4</intersection>
<intersection>62 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>57,-34.5,57,-33</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<intersection>-34.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-33.5,50,-27</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<connection>
<GID>139</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>52,-27,56,-27</points>
<connection>
<GID>142</GID>
<name>OUT</name></connection>
<connection>
<GID>140</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>51,-21,51,-21</points>
<connection>
<GID>140</GID>
<name>OUT</name></connection>
<connection>
<GID>149</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-27,61,-21</points>
<connection>
<GID>141</GID>
<name>OUT</name></connection>
<connection>
<GID>150</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-46,44.5,-19</points>
<intersection>-46 2</intersection>
<intersection>-19 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>38,-46,38,-45</points>
<connection>
<GID>130</GID>
<name>N_in0</name></connection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>38,-46,44.5,-46</points>
<intersection>38 1</intersection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>44.5,-19,51,-19</points>
<connection>
<GID>149</GID>
<name>N_in1</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-46,62,-45</points>
<connection>
<GID>145</GID>
<name>N_in0</name></connection>
<intersection>-46 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>68.5,-46,68.5,-19</points>
<intersection>-46 2</intersection>
<intersection>-19 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>62,-46,68.5,-46</points>
<intersection>62 0</intersection>
<intersection>68.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>68.5,-19,75,-19</points>
<connection>
<GID>98</GID>
<name>N_in1</name></connection>
<intersection>68.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86,-72,97,-72</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>97 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>97,-77,97,-45</points>
<connection>
<GID>113</GID>
<name>N_in0</name></connection>
<connection>
<GID>154</GID>
<name>N_in3</name></connection>
<intersection>-72 1</intersection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94,-77,94,-49.5</points>
<connection>
<GID>155</GID>
<name>N_in3</name></connection>
<intersection>-70 1</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86,-70,94,-70</points>
<connection>
<GID>153</GID>
<name>OUT_1</name></connection>
<intersection>94 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73,-49.5,94,-49.5</points>
<intersection>73 3</intersection>
<intersection>94 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>73,-49.5,73,-45</points>
<connection>
<GID>90</GID>
<name>N_in0</name></connection>
<intersection>-49.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-77,91,-55.5</points>
<connection>
<GID>156</GID>
<name>N_in3</name></connection>
<intersection>-68 5</intersection>
<intersection>-55.5 7</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>86,-68,91,-68</points>
<connection>
<GID>153</GID>
<name>OUT_2</name></connection>
<intersection>91 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>49,-55.5,91,-55.5</points>
<intersection>49 8</intersection>
<intersection>91 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>49,-55.5,49,-45</points>
<connection>
<GID>143</GID>
<name>N_in0</name></connection>
<intersection>-55.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-77,88,-59.5</points>
<connection>
<GID>157</GID>
<name>N_in3</name></connection>
<intersection>-66 9</intersection>
<intersection>-59.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>25,-59.5,88,-59.5</points>
<intersection>25 7</intersection>
<intersection>88 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>25,-59.5,25,-45</points>
<connection>
<GID>128</GID>
<name>N_in0</name></connection>
<intersection>-59.5 6</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>86,-66,88,-66</points>
<connection>
<GID>153</GID>
<name>OUT_3</name></connection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,-29,109,-9</points>
<connection>
<GID>160</GID>
<name>N_in2</name></connection>
<connection>
<GID>120</GID>
<name>N_in1</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109,-15,118.5,-15</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>109 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-19,85,-14</points>
<connection>
<GID>101</GID>
<name>N_in1</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-14,118.5,-14</points>
<connection>
<GID>159</GID>
<name>IN_1</name></connection>
<intersection>85 0</intersection>
<intersection>106 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>106,-14,106,-8</points>
<connection>
<GID>161</GID>
<name>N_in2</name></connection>
<intersection>-14 1</intersection>
<intersection>-8 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>105,-8,106,-8</points>
<connection>
<GID>161</GID>
<name>N_in0</name></connection>
<intersection>106 2</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-19,61,-13</points>
<connection>
<GID>150</GID>
<name>N_in1</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-13,118.5,-13</points>
<connection>
<GID>159</GID>
<name>IN_2</name></connection>
<intersection>61 0</intersection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-13,103,-9</points>
<connection>
<GID>162</GID>
<name>N_in2</name></connection>
<intersection>-13 1</intersection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-19,37,-12</points>
<connection>
<GID>135</GID>
<name>N_in1</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-12,118.5,-12</points>
<connection>
<GID>159</GID>
<name>IN_3</name></connection>
<intersection>37 0</intersection>
<intersection>100 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>100,-12,100,-9</points>
<connection>
<GID>163</GID>
<name>N_in2</name></connection>
<intersection>-12 1</intersection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-19,27,-11</points>
<connection>
<GID>134</GID>
<name>N_in1</name></connection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27,-11,95,-11</points>
<intersection>27 0</intersection>
<intersection>95 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>95,-11,95,-9</points>
<connection>
<GID>165</GID>
<name>N_in2</name></connection>
<intersection>-11 2</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-69.4231,23.183,108.608,-68.7365</PageViewport>
<gate>
<ID>2</ID>
<type>AA_FULLADDER_1BIT</type>
<position>28,-19.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_B_0</ID>15 </input>
<output>
<ID>OUT_0</ID>23 </output>
<input>
<ID>carry_in</ID>7 </input>
<output>
<ID>carry_out</ID>11 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_FULLADDER_1BIT</type>
<position>39.5,-19.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_B_0</ID>14 </input>
<output>
<ID>OUT_0</ID>22 </output>
<input>
<ID>carry_in</ID>8 </input>
<output>
<ID>carry_out</ID>7 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_FULLADDER_1BIT</type>
<position>51,-19.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_B_0</ID>13 </input>
<output>
<ID>OUT_0</ID>21 </output>
<input>
<ID>carry_in</ID>9 </input>
<output>
<ID>carry_out</ID>8 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_FULLADDER_1BIT</type>
<position>62.5,-19.5</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_B_0</ID>12 </input>
<output>
<ID>OUT_0</ID>20 </output>
<input>
<ID>carry_in</ID>10 </input>
<output>
<ID>carry_out</ID>9 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7</ID>
<type>DD_KEYPAD_HEX</type>
<position>17.5,4.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<output>
<ID>OUT_1</ID>13 </output>
<output>
<ID>OUT_2</ID>14 </output>
<output>
<ID>OUT_3</ID>15 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>11</ID>
<type>DD_KEYPAD_HEX</type>
<position>17.5,-9</position>
<output>
<ID>OUT_0</ID>16 </output>
<output>
<ID>OUT_1</ID>17 </output>
<output>
<ID>OUT_2</ID>18 </output>
<output>
<ID>OUT_3</ID>19 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>FF_GND</type>
<position>68,-20.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>19.5,-19.5</position>
<input>
<ID>N_in1</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>14,-19</position>
<gparam>LABEL_TEXT Overflow</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>75,-28</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<input>
<ID>IN_2</ID>22 </input>
<input>
<ID>IN_3</ID>23 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>12,4.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>12,-8.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>74.5,-22.5</position>
<gparam>LABEL_TEXT SUM</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,-19.5,35.5,-19.5</points>
<connection>
<GID>2</GID>
<name>carry_in</name></connection>
<connection>
<GID>3</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43.5,-19.5,47,-19.5</points>
<connection>
<GID>3</GID>
<name>carry_in</name></connection>
<connection>
<GID>4</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-19.5,58.5,-19.5</points>
<connection>
<GID>4</GID>
<name>carry_in</name></connection>
<connection>
<GID>5</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>66.5,-19.5,68,-19.5</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<connection>
<GID>5</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-19.5,24,-19.5</points>
<connection>
<GID>2</GID>
<name>carry_out</name></connection>
<connection>
<GID>18</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-16.5,61.5,1.5</points>
<connection>
<GID>5</GID>
<name>IN_B_0</name></connection>
<intersection>1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,1.5,61.5,1.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-16.5,50,3.5</points>
<connection>
<GID>4</GID>
<name>IN_B_0</name></connection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,3.5,50,3.5</points>
<connection>
<GID>7</GID>
<name>OUT_1</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-16.5,38.5,5.5</points>
<connection>
<GID>3</GID>
<name>IN_B_0</name></connection>
<intersection>5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,5.5,38.5,5.5</points>
<connection>
<GID>7</GID>
<name>OUT_2</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-16.5,27,7.5</points>
<connection>
<GID>2</GID>
<name>IN_B_0</name></connection>
<intersection>7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,7.5,27,7.5</points>
<connection>
<GID>7</GID>
<name>OUT_3</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-16.5,63.5,-12</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-12,63.5,-12</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-16.5,52,-10</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-10,52,-10</points>
<connection>
<GID>11</GID>
<name>OUT_1</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-16.5,40.5,-8</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-8,40.5,-8</points>
<connection>
<GID>11</GID>
<name>OUT_2</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-16.5,29,-6</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-6,29,-6</points>
<connection>
<GID>11</GID>
<name>OUT_3</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-29,62.5,-22.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-29,72,-29</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-28,51,-22.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-28,72,-28</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-27,72,-27</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<intersection>39.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>39.5,-27,39.5,-22.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>-27 1</intersection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-26,28,-22.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-26,72,-26</points>
<connection>
<GID>22</GID>
<name>IN_3</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>34.9113,-12.4986,212.943,-104.418</PageViewport>
<gate>
<ID>27</ID>
<type>AA_FULLADDER_1BIT</type>
<position>86.5,-66.5</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_B_0</ID>32 </input>
<output>
<ID>OUT_0</ID>40 </output>
<input>
<ID>carry_in</ID>24 </input>
<output>
<ID>carry_out</ID>28 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_FULLADDER_1BIT</type>
<position>98,-66.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_B_0</ID>31 </input>
<output>
<ID>OUT_0</ID>39 </output>
<input>
<ID>carry_in</ID>25 </input>
<output>
<ID>carry_out</ID>24 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_FULLADDER_1BIT</type>
<position>109.5,-66.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_B_0</ID>30 </input>
<output>
<ID>OUT_0</ID>38 </output>
<input>
<ID>carry_in</ID>26 </input>
<output>
<ID>carry_out</ID>25 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_FULLADDER_1BIT</type>
<position>121,-66.5</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_B_0</ID>29 </input>
<output>
<ID>OUT_0</ID>37 </output>
<input>
<ID>carry_in</ID>59 </input>
<output>
<ID>carry_out</ID>26 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>31</ID>
<type>DD_KEYPAD_HEX</type>
<position>67.5,-34.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<output>
<ID>OUT_1</ID>30 </output>
<output>
<ID>OUT_2</ID>31 </output>
<output>
<ID>OUT_3</ID>32 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>DD_KEYPAD_HEX</type>
<position>67.5,-51.5</position>
<output>
<ID>OUT_0</ID>41 </output>
<output>
<ID>OUT_1</ID>44 </output>
<output>
<ID>OUT_2</ID>47 </output>
<output>
<ID>OUT_3</ID>51 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>78,-66.5</position>
<input>
<ID>N_in1</ID>28 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>72.5,-66</position>
<gparam>LABEL_TEXT Overflow</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>133.5,-75</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>39 </input>
<input>
<ID>IN_3</ID>40 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>62,-34.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>62,-51.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>133,-69.5</position>
<gparam>LABEL_TEXT X+Y/X-Y</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AI_XOR2</type>
<position>79.5,-48.5</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AI_XOR2</type>
<position>79.5,-53.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>AI_XOR2</type>
<position>79.5,-58.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AI_XOR2</type>
<position>79.5,-43.5</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>66,-62</position>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>63,-61.5</position>
<gparam>LABEL_TEXT +/-</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>90.5,-66.5,94,-66.5</points>
<connection>
<GID>27</GID>
<name>carry_in</name></connection>
<connection>
<GID>28</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>102,-66.5,105.5,-66.5</points>
<connection>
<GID>28</GID>
<name>carry_in</name></connection>
<connection>
<GID>29</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>113.5,-66.5,117,-66.5</points>
<connection>
<GID>29</GID>
<name>carry_in</name></connection>
<connection>
<GID>30</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79,-66.5,82.5,-66.5</points>
<connection>
<GID>34</GID>
<name>N_in1</name></connection>
<connection>
<GID>27</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-63.5,120,-37.5</points>
<connection>
<GID>30</GID>
<name>IN_B_0</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-37.5,120,-37.5</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-63.5,108.5,-35.5</points>
<connection>
<GID>29</GID>
<name>IN_B_0</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-35.5,108.5,-35.5</points>
<connection>
<GID>31</GID>
<name>OUT_1</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-63.5,97,-33.5</points>
<connection>
<GID>28</GID>
<name>IN_B_0</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-33.5,97,-33.5</points>
<connection>
<GID>31</GID>
<name>OUT_2</name></connection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-63.5,85.5,-31.5</points>
<connection>
<GID>27</GID>
<name>IN_B_0</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-31.5,85.5,-31.5</points>
<connection>
<GID>31</GID>
<name>OUT_3</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-76,121,-69.5</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>-76 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-76,130.5,-76</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-75,109.5,-69.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,-75,130.5,-75</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-74,130.5,-74</points>
<connection>
<GID>36</GID>
<name>IN_2</name></connection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-74,98,-69.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>-74 1</intersection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-73,86.5,-69.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,-73,130.5,-73</points>
<connection>
<GID>36</GID>
<name>IN_3</name></connection>
<intersection>86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-57.5,73,-54.5</points>
<intersection>-57.5 2</intersection>
<intersection>-54.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>73,-57.5,76.5,-57.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>72.5,-54.5,73,-54.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72.5,-52.5,76.5,-52.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<connection>
<GID>32</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-50.5,73.5,-47.5</points>
<intersection>-50.5 1</intersection>
<intersection>-47.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-50.5,73.5,-50.5</points>
<connection>
<GID>32</GID>
<name>OUT_2</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-47.5,76.5,-47.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-48.5,72.5,-42.5</points>
<connection>
<GID>32</GID>
<name>OUT_3</name></connection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>72.5,-42.5,76.5,-42.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-63.5,122,-58.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-58.5,122,-58.5</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>122 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-63.5,110.5,-53.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-53.5,110.5,-53.5</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-63.5,99,-48.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-48.5,99,-48.5</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-63.5,87.5,-43.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-43.5,87.5,-43.5</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-62,74.5,-44.5</points>
<intersection>-62 1</intersection>
<intersection>-59.5 8</intersection>
<intersection>-54.5 4</intersection>
<intersection>-49.5 3</intersection>
<intersection>-44.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-62,125,-62</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>74.5 0</intersection>
<intersection>125 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74.5,-44.5,76.5,-44.5</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>74.5,-49.5,76.5,-49.5</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>74.5,-54.5,76.5,-54.5</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>125,-66.5,125,-62</points>
<connection>
<GID>30</GID>
<name>carry_in</name></connection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>74.5,-59.5,76.5,-59.5</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-77.0226,30.6543,160.353,-91.9051</PageViewport>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>23.5,-12</position>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_TOGGLE</type>
<position>23.5,-20</position>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_AND2</type>
<position>38,-13</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>19.5,-11.5</position>
<gparam>LABEL_TEXT IP</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>20,-19.5</position>
<gparam>LABEL_TEXT M</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>53.5,-13</position>
<input>
<ID>N_in0</ID>63 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>56.5,-12.5</position>
<gparam>LABEL_TEXT N</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>39,-3</position>
<gparam>LABEL_TEXT 32x</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AE_SMALL_INVERTER</type>
<position>-175,18.5</position>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_INVERTER</type>
<position>38,-20</position>
<input>
<ID>IN_0</ID>61 </input>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>68</ID>
<type>AE_OR2</type>
<position>46,-19</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>GA_LED</type>
<position>53.5,-19</position>
<input>
<ID>N_in0</ID>93 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>56.5,-18.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-12,35,-12</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<connection>
<GID>53</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-20,30.5,-14</points>
<intersection>-20 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-20,35,-20</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-14,35,-14</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-13,52.5,-13</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<connection>
<GID>59</GID>
<name>N_in0</name></connection>
<intersection>43 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>43,-18,43,-13</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>-13 1</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-20,43,-20</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,-19,52.5,-19</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<connection>
<GID>70</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>-1.9031e-006,8.32477,316.5,-155.088</PageViewport></page 4>
<page 5>
<PageViewport>-1.9031e-006,8.32477,316.5,-155.088</PageViewport></page 5>
<page 6>
<PageViewport>-1.9031e-006,8.32477,316.5,-155.088</PageViewport></page 6>
<page 7>
<PageViewport>-1.9031e-006,8.32477,316.5,-155.088</PageViewport></page 7>
<page 8>
<PageViewport>-1.9031e-006,8.32477,316.5,-155.088</PageViewport></page 8>
<page 9>
<PageViewport>-1.9031e-006,8.32477,316.5,-155.088</PageViewport></page 9></circuit>