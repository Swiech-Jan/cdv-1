<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>1.63402,2.88289,51.2465,-31.1484</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>10,-0.5</position>
<gparam>LABEL_TEXT Y = !ABC + A!C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AE_OR2</type>
<position>36,-19.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND3</type>
<position>26.5,-16.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>4 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_AND2</type>
<position>26.5,-26.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>6.5,-3.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>4.5,-3</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>6.5,-7</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>4.5,-6.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>6.5,-10.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>4.5,-10</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_INVERTER</type>
<position>18.5,-13</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>20</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>44,-18.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_INVERTER</type>
<position>15,-27.5</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-13,13.5,-3.5</points>
<intersection>-13 1</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13.5,-13,15.5,-13</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>13.5 0</intersection>
<intersection>15.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-3.5,13.5,-3.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>13.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15.5,-25.5,15.5,-13</points>
<intersection>-25.5 4</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>15.5,-25.5,23.5,-25.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-14.5,23.5,-14.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>21.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>21.5,-14.5,21.5,-13</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-16.5,12,-7</points>
<intersection>-16.5 1</intersection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-16.5,23.5,-16.5</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-7,12,-7</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>12 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-18.5,10.5,-10.5</points>
<intersection>-18.5 1</intersection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-18.5,23.5,-18.5</points>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<intersection>10.5 0</intersection>
<intersection>12 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-10.5,10.5,-10.5</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>10.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>12,-27.5,12,-18.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-18.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-18.5,31,-16.5</points>
<intersection>-18.5 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-18.5,33,-18.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-16.5,31,-16.5</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-19.5,41,-19.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,-27.5,23.5,-27.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-26.5,31,-20.5</points>
<intersection>-26.5 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-20.5,33,-20.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-26.5,31,-26.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-2.475,1.45,63.675,-43.925</PageViewport>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>4.5,-0.5</position>
<gparam>LABEL_TEXT Y = !AB + !ACD</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>2,-4.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>-0.5,-4</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>2,-7.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>-0.5,-7</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_TOGGLE</type>
<position>2,-10.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>-0.5,-10</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>2,-13.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>-0.5,-13</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AE_OR2</type>
<position>39,-22</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_AND2</type>
<position>28.5,-18.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_AND3</type>
<position>28.5,-25.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>12 </input>
<input>
<ID>IN_2</ID>13 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_INVERTER</type>
<position>17.5,-15.5</position>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>44</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>46.5,-21</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-15.5,13,-4.5</points>
<intersection>-15.5 1</intersection>
<intersection>-4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-15.5,14.5,-15.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4,-4.5,13,-4.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>13 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-15.5,23,-15.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>23 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>23,-23.5,23,-15.5</points>
<intersection>-23.5 9</intersection>
<intersection>-17.5 10</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>23,-23.5,25.5,-23.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>23 7</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>23,-17.5,25.5,-17.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>23 7</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-19.5,11,-7.5</points>
<intersection>-19.5 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-7.5,11,-7.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-19.5,25.5,-19.5</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-25.5,9,-10.5</points>
<intersection>-25.5 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-10.5,9,-10.5</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9,-25.5,25.5,-25.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-27.5,7,-13.5</points>
<intersection>-27.5 2</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-13.5,7,-13.5</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>7 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7,-27.5,25.5,-27.5</points>
<connection>
<GID>40</GID>
<name>IN_2</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-21,33.5,-18.5</points>
<intersection>-21 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-21,36,-21</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-18.5,33.5,-18.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-25.5,33.5,-23</points>
<intersection>-25.5 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-23,36,-23</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-25.5,33.5,-25.5</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42,-22,43.5,-22</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<connection>
<GID>36</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-4.725,1.45,61.425,-43.925</PageViewport>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>5.5,-0.5</position>
<gparam>LABEL_TEXT Y = !A(B+C) (B+D)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_AND3</type>
<position>31.5,-19</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>22 </input>
<input>
<ID>IN_2</ID>23 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>50</ID>
<type>AE_OR2</type>
<position>16,-17</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>AE_OR2</type>
<position>16,-25</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_TOGGLE</type>
<position>2,-4.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>-0.5,-4</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>2,-7</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>-0.5,-6.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_TOGGLE</type>
<position>2,-9.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>-0.5,-9</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_TOGGLE</type>
<position>2,-12</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>-0.5,-11.5</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_INVERTER</type>
<position>16,-4.5</position>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>66</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>40.5,-18</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-4.5,13,-4.5</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<connection>
<GID>64</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-17,23.5,-4.5</points>
<intersection>-17 1</intersection>
<intersection>-4.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-17,28.5,-17</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>19,-4.5,23.5,-4.5</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-16,11,-7</points>
<intersection>-16 1</intersection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,-16,13,-16</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>11 0</intersection>
<intersection>12 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4,-7,11,-7</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>11 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>12,-24,12,-16</points>
<intersection>-24 4</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>12,-24,13,-24</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>12 3</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-18,9,-9.5</points>
<intersection>-18 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-18,13,-18</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4,-9.5,9,-9.5</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-26,7,-12</points>
<intersection>-26 2</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-12,7,-12</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<intersection>7 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7,-26,13,-26</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-19,21.5,-17</points>
<intersection>-19 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-19,28.5,-19</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19,-17,21.5,-17</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-25,23.5,-21</points>
<intersection>-25 2</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-21,28.5,-21</points>
<connection>
<GID>48</GID>
<name>IN_2</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19,-25,23.5,-25</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-19,37.5,-19</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<connection>
<GID>48</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,0,88.2,-60.5</PageViewport>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>14.5,-1.5</position>
<gparam>LABEL_TEXT Uklad sumujacy (funkcja S oraz C)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_TOGGLE</type>
<position>3.5,-6.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>3.5,-4</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AA_TOGGLE</type>
<position>13,-6.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>13,-4</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AA_TOGGLE</type>
<position>23.5,-6.5</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>23.5,-4</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AE_OR2</type>
<position>55.5,-17.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>AE_OR3</type>
<position>56,-37.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<input>
<ID>IN_2</ID>36 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>82</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>64.5,-16.5</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>83</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>64.5,-36.5</position>
<input>
<ID>IN_0</ID>37 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_AND2</type>
<position>44.5,-12.5</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_AND2</type>
<position>46.5,-20</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>88</ID>
<type>AA_AND2</type>
<position>45,-31</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>AA_AND2</type>
<position>45,-37.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_AND2</type>
<position>45,-43.5</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>AO_XNOR2</type>
<position>36,-10.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_INVERTER</type>
<position>38.5,-24</position>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>96</ID>
<type>AI_XOR2</type>
<position>38.5,-18.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_LABEL</type>
<position>64.5,-11</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>AA_LABEL</type>
<position>64.5,-31</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-9.5,10.5,-6.5</points>
<intersection>-9.5 1</intersection>
<intersection>-6.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-9.5,33,-9.5</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>10.5 0</intersection>
<intersection>17.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5.5,-6.5,10.5,-6.5</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<intersection>10.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>17.5,-17.5,17.5,-9.5</points>
<intersection>-17.5 4</intersection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>17.5,-17.5,35.5,-17.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>17.5 3</intersection>
<intersection>22.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>22.5,-30,22.5,-17.5</points>
<intersection>-30 6</intersection>
<intersection>-17.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>22.5,-30,42,-30</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>22.5 5</intersection>
<intersection>33 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>33,-36.5,33,-30</points>
<intersection>-36.5 8</intersection>
<intersection>-30 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>33,-36.5,42,-36.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>33 7</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-11.5,20.5,-6.5</points>
<intersection>-11.5 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-6.5,20.5,-6.5</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20.5,-11.5,33,-11.5</points>
<connection>
<GID>92</GID>
<name>IN_1</name></connection>
<intersection>20.5 0</intersection>
<intersection>24 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24,-19.5,24,-11.5</points>
<intersection>-19.5 4</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>24,-19.5,35.5,-19.5</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>24 3</intersection>
<intersection>29 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>29,-38.5,29,-19.5</points>
<intersection>-38.5 6</intersection>
<intersection>-19.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>29,-38.5,42,-38.5</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<intersection>29 5</intersection>
<intersection>33 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>33,-42.5,33,-38.5</points>
<intersection>-42.5 8</intersection>
<intersection>-38.5 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>33,-42.5,42,-42.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>33 7</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-10.5,41.5,-10.5</points>
<connection>
<GID>92</GID>
<name>OUT</name></connection>
<intersection>41.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>41.5,-11.5,41.5,-10.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>-10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-13.5,29,-6.5</points>
<intersection>-13.5 1</intersection>
<intersection>-6.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-13.5,41.5,-13.5</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection>
<intersection>33 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-6.5,29,-6.5</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33,-24,33,-13.5</points>
<intersection>-24 4</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>33,-24,35.5,-24</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>33 3</intersection>
<intersection>35.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>35.5,-32,35.5,-24</points>
<intersection>-32 6</intersection>
<intersection>-24 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>35.5,-32,42,-32</points>
<connection>
<GID>88</GID>
<name>IN_1</name></connection>
<intersection>35.5 5</intersection>
<intersection>38 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>38,-44.5,38,-32</points>
<intersection>-44.5 8</intersection>
<intersection>-32 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>38,-44.5,42,-44.5</points>
<connection>
<GID>90</GID>
<name>IN_1</name></connection>
<intersection>38 7</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-16.5,50,-12.5</points>
<intersection>-16.5 1</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-16.5,52.5,-16.5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47.5,-12.5,50,-12.5</points>
<connection>
<GID>85</GID>
<name>OUT</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41.5,-24,43.5,-24</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>43.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>43.5,-24,43.5,-21</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<intersection>-24 1</intersection></vsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-19,42.5,-18.5</points>
<intersection>-19 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-19,43.5,-19</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-18.5,42.5,-18.5</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-20,51,-18.5</points>
<intersection>-20 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-18.5,52.5,-18.5</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-20,51,-20</points>
<connection>
<GID>86</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-17.5,61.5,-17.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<connection>
<GID>78</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-35.5,49.5,-31</points>
<intersection>-35.5 1</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-35.5,53,-35.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-31,49.5,-31</points>
<connection>
<GID>88</GID>
<name>OUT</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-37.5,53,-37.5</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<connection>
<GID>89</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-43.5,49.5,-39.5</points>
<intersection>-43.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-39.5,53,-39.5</points>
<connection>
<GID>80</GID>
<name>IN_2</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-43.5,49.5,-43.5</points>
<connection>
<GID>90</GID>
<name>OUT</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59,-37.5,61.5,-37.5</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<connection>
<GID>83</GID>
<name>IN_0</name></connection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>-8.53137,6.93914,57.6186,-38.4359</PageViewport>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>-2.5,5</position>
<gparam>LABEL_TEXT Polsumator</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>AA_TOGGLE</type>
<position>-3.5,1</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>-6,1.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_TOGGLE</type>
<position>-3.5,-2.5</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>-6,-2</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>AE_OR2</type>
<position>28,-14.5</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_AND2</type>
<position>19.5,-9.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_AND2</type>
<position>19.5,-20</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_INVERTER</type>
<position>10,-12.5</position>
<input>
<ID>IN_0</ID>40 </input>
<output>
<ID>OUT_0</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>117</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>36.5,-12.5</position>
<input>
<ID>IN_0</ID>41 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>36.5,-7</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>119</ID>
<type>AA_INVERTER</type>
<position>10,-17.5</position>
<input>
<ID>IN_0</ID>38 </input>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_AND2</type>
<position>27.5,-27.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>122</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>36.5,-26.5</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_LABEL</type>
<position>36.5,-21</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-8.5,3.5,1</points>
<intersection>-8.5 2</intersection>
<intersection>1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1.5,1,3.5,1</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<intersection>3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3.5,-8.5,16.5,-8.5</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>3.5 0</intersection>
<intersection>5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>5,-17.5,5,-8.5</points>
<intersection>-17.5 4</intersection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>5,-17.5,7,-17.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>5 3</intersection>
<intersection>7 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>7,-26.5,7,-17.5</points>
<intersection>-26.5 6</intersection>
<intersection>-17.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>7,-26.5,24.5,-26.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>7 5</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-12.5,14.5,-10.5</points>
<intersection>-12.5 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-10.5,16.5,-10.5</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-12.5,14.5,-12.5</points>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-0.5,-12.5,-0.5,-2.5</points>
<intersection>-12.5 2</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1.5,-2.5,-0.5,-2.5</points>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection>
<intersection>-0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-0.5,-12.5,7,-12.5</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>-0.5 0</intersection>
<intersection>1.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1.5,-21,1.5,-12.5</points>
<intersection>-21 4</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>1.5,-21,16.5,-21</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<intersection>1.5 3</intersection>
<intersection>13.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>13.5,-28.5,13.5,-21</points>
<intersection>-28.5 6</intersection>
<intersection>-21 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>13.5,-28.5,24.5,-28.5</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>13.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-14.5,33.5,-14.5</points>
<connection>
<GID>110</GID>
<name>OUT</name></connection>
<intersection>33.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>33.5,-14.5,33.5,-13.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>-14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-13.5,24.5,-9.5</points>
<intersection>-13.5 3</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-9.5,24.5,-9.5</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24.5,-13.5,25,-13.5</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-19,14.5,-17.5</points>
<intersection>-19 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-19,16.5,-19</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-17.5,14.5,-17.5</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-20,23.5,-15.5</points>
<intersection>-20 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-15.5,25,-15.5</points>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-20,23.5,-20</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-27.5,33.5,-27.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<connection>
<GID>121</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>-2.475,1.45,63.675,-43.925</PageViewport>
<gate>
<ID>125</ID>
<type>AA_TOGGLE</type>
<position>1,-3</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>-1,-2.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>3.5,0</position>
<gparam>LABEL_TEXT Polsumator</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>AA_TOGGLE</type>
<position>1,-6</position>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_LABEL</type>
<position>-1,-5.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AI_XOR2</type>
<position>13.5,-9.5</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>21.5,-8.5</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>135</ID>
<type>AA_LABEL</type>
<position>21.5,-3</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>137</ID>
<type>AA_AND2</type>
<position>13.5,-18</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>21.5,-18.5</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>139</ID>
<type>AA_LABEL</type>
<position>21.5,-13</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-8.5,8,-3</points>
<intersection>-8.5 1</intersection>
<intersection>-3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,-8.5,10.5,-8.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection>
<intersection>9 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3,-3,8,-3</points>
<connection>
<GID>125</GID>
<name>OUT_0</name></connection>
<intersection>8 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>9,-17,9,-8.5</points>
<intersection>-17 4</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>9,-17,10.5,-17</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>9 3</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-10.5,6.5,-6</points>
<intersection>-10.5 1</intersection>
<intersection>-6 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-10.5,10.5,-10.5</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>6.5 0</intersection>
<intersection>7.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3,-6,6.5,-6</points>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection>
<intersection>6.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>7.5,-19,7.5,-10.5</points>
<intersection>-19 4</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>7.5,-19,10.5,-19</points>
<connection>
<GID>137</GID>
<name>IN_1</name></connection>
<intersection>7.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-9.5,18.5,-9.5</points>
<connection>
<GID>132</GID>
<name>OUT</name></connection>
<connection>
<GID>134</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-19.5,17.5,-18</points>
<intersection>-19.5 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-19.5,18.5,-19.5</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-18,17.5,-18</points>
<connection>
<GID>137</GID>
<name>OUT</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>0,0,88.2,-60.5</PageViewport>
<gate>
<ID>141</ID>
<type>AA_LABEL</type>
<position>5,-2</position>
<gparam>LABEL_TEXT Sumator</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>AE_OR4</type>
<position>30,-26</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>51 </input>
<input>
<ID>IN_2</ID>52 </input>
<input>
<ID>IN_3</ID>53 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_AND3</type>
<position>12.5,-9.5</position>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_LABEL</type>
<position>8,-7</position>
<gparam>LABEL_TEXT !A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>AA_LABEL</type>
<position>8,-9</position>
<gparam>LABEL_TEXT !B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>AA_LABEL</type>
<position>7,-11</position>
<gparam>LABEL_TEXT C (IN)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>AA_AND3</type>
<position>12.5,-18</position>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_LABEL</type>
<position>8,-15.5</position>
<gparam>LABEL_TEXT !A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>AA_LABEL</type>
<position>8,-17.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>AA_LABEL</type>
<position>6.5,-19.5</position>
<gparam>LABEL_TEXT !C (IN)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>AA_AND3</type>
<position>12.5,-27</position>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_LABEL</type>
<position>8,-24.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>AA_LABEL</type>
<position>8,-26.5</position>
<gparam>LABEL_TEXT !B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>AA_LABEL</type>
<position>6.5,-28.5</position>
<gparam>LABEL_TEXT !C (IN)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>AA_AND3</type>
<position>12.5,-35.5</position>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_LABEL</type>
<position>8,-33</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>AA_LABEL</type>
<position>8,-35</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>AA_LABEL</type>
<position>6.5,-37</position>
<gparam>LABEL_TEXT C (IN)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>AA_LABEL</type>
<position>35.5,-25.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>AE_OR3</type>
<position>65.5,-28</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>55 </input>
<input>
<ID>IN_2</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>168</ID>
<type>AA_AND2</type>
<position>53.5,-21.5</position>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>169</ID>
<type>AA_LABEL</type>
<position>48.5,-20</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AA_LABEL</type>
<position>48.5,-22</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>AA_AND2</type>
<position>53.5,-27</position>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_LABEL</type>
<position>48.5,-25.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>AA_LABEL</type>
<position>47.5,-27.5</position>
<gparam>LABEL_TEXT C (IN)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>AA_AND2</type>
<position>53.5,-32.5</position>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>175</ID>
<type>AA_LABEL</type>
<position>48.5,-31</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>176</ID>
<type>AA_LABEL</type>
<position>47.5,-33</position>
<gparam>LABEL_TEXT C (IN)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-23,23.5,-9.5</points>
<intersection>-23 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-23,27,-23</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,-9.5,23.5,-9.5</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-25,22,-18</points>
<intersection>-25 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-25,27,-25</points>
<connection>
<GID>143</GID>
<name>IN_1</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,-18,22,-18</points>
<connection>
<GID>152</GID>
<name>OUT</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15.5,-27,27,-27</points>
<connection>
<GID>156</GID>
<name>OUT</name></connection>
<connection>
<GID>143</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-35.5,23.5,-29</points>
<intersection>-35.5 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-29,27,-29</points>
<connection>
<GID>143</GID>
<name>IN_3</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,-35.5,23.5,-35.5</points>
<connection>
<GID>160</GID>
<name>OUT</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-26,59.5,-21.5</points>
<intersection>-26 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,-26,62.5,-26</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-21.5,59.5,-21.5</points>
<connection>
<GID>168</GID>
<name>OUT</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-28,59.5,-27</points>
<intersection>-28 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,-28,62.5,-28</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-27,59.5,-27</points>
<connection>
<GID>171</GID>
<name>OUT</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-32.5,59.5,-30</points>
<intersection>-32.5 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,-30,62.5,-30</points>
<connection>
<GID>166</GID>
<name>IN_2</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-32.5,59.5,-32.5</points>
<connection>
<GID>174</GID>
<name>OUT</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire></page 6>
<page 7>
<PageViewport>0,0,88.2,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,88.2,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,88.2,-60.5</PageViewport></page 9></circuit>